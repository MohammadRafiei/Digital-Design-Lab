module dec4to16(A,C,B,D,y);
input A,C,B,D;
output [15:0] y;
wire A0,B0,C0,D0, f1,f2,f3,f4;
not(A0,A);
not(B0,B);
not(C0,C);
not(D0,D);
// and(f1,E,A0,B0);
// and(f2,E.A0,B);
// and(f3,E,A0,B0);
// and(f4,E,A,B);
and(y[0],f1,C0,D0);
and(y[1],f1,C0,D);
and(y[2],f1,C,D0);
and(y[3],f1,C,D);
and(y[4],f2,C0,D0);
and(y[5],f2,C0,D);
and(y[6],f2,C,D0);
and(y[7],f2,C,D);
and(y[8],f3,C0,D0);
and(y[9],f3,C0,D);
and(y[10],f3,C,D0);
and(y[11],f3,C,D);
and(y[12],f4,C0,D0);
and(y[13],f4,C0,D);
and(y[14],f4,C,D0);
and(y[15],f4,C,D);
endmodule