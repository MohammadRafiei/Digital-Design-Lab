module add(input1,input2,output3);
input  [31:0] input1, input2;
output [31:0] out;

	assign output3 = input1 + input2;
endmodule